architecture behavioral of ent is
begin

    signal_name <= 	expression_1 when condition_1 else
                    expression_2 when condition_2 else
                    expression_3 ;

end behavioral ; -- arch
