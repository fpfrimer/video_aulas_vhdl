
-- Exemplo de rótulo, utilizado para facilitar 
-- o entendimento dos códigos

nome_rotulo: block
    -- Definiçâo de sinais
begin
    -- Comandos concorrentes
    -- Comandos concorrentes
end block nome_rotulo;